// axi-constants.svh
`include "axi_constants.svh"

// axi-base
`include "IfAxi.sv"
`include "TrAxi.sv"

// axi-channel
`include "AxiMstrChnAw.sv"
`include "AxiMstrChnW.sv"
`include "AxiMstrChnB.sv"
`include "AxiMstrChnAr.sv"
`include "AxiMstrChnR.sv"

// axi-agent
`include "AxiMstrSqr.sv"
`include "AxiMstrAgtWr.sv"
`include "AxiMstrAgtRd.sv"

// axi-env
`include "AxiSlvRef.sv"
`include "AxiSlvScb.sv"
`include "AxiMstrVirSqrWr.sv"
`include "AxiMstrEnv.sv"

// axi-seq
`include "AxiMstrSeqWr.sv"
`include "AxiMstrSeqRd.sv"




